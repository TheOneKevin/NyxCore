module hs32_lsu (
    input wire clk,
    input wire reset
);
    
endmodule