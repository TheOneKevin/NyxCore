`default_nettype none

`include "rtl/include/utils.svh"
`include "rtl/include/types.svh"
`include "rtl/hs32_lcu.sv"
`include "rtl/hs32_adder.sv"
`include "rtl/hs32_alu.sv"
`include "rtl/hs32_primitives.sv"
`include "rtl/hs32_regfile4r1w.sv"
`include "rtl/hs32_decode1.sv"
`include "rtl/hs32_decode2.sv"
`include "rtl/hs32_execute.sv"
`include "rtl/hs32_pipeline.sv"
