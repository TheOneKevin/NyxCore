`include "primitives/skid_buffer.svh"
`include "primitives/shift_right.svh"
`include "primitives/mux2to1.svh"
`include "primitives/mux4to1.svh"