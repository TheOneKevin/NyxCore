module sram_wrapper #(
    parameter ADDR_WIDTH = 10,
    parameter NUM_RP     = 1,
    parameter NUM_WP     = 2
) (
    ports
);
    
endmodule